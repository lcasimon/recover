magic
tech sky130A
timestamp 1694812110
<< pwell >>
rect -123 -180 123 180
<< nmos >>
rect -25 -75 25 75
<< ndiff >>
rect -54 69 -25 75
rect -54 -69 -48 69
rect -31 -69 -25 69
rect -54 -75 -25 -69
rect 25 69 54 75
rect 25 -69 31 69
rect 48 -69 54 69
rect 25 -75 54 -69
<< ndiffc >>
rect -48 -69 -31 69
rect 31 -69 48 69
<< psubdiff >>
rect -105 145 -57 162
rect 57 145 105 162
rect -105 114 -88 145
rect 88 114 105 145
rect -105 -145 -88 -114
rect 88 -145 105 -114
rect -105 -162 -57 -145
rect 57 -162 105 -145
<< psubdiffcont >>
rect -57 145 57 162
rect -105 -114 -88 114
rect 88 -114 105 114
rect -57 -162 57 -145
<< poly >>
rect -25 111 25 119
rect -25 94 -17 111
rect 17 94 25 111
rect -25 75 25 94
rect -25 -94 25 -75
rect -25 -111 -17 -94
rect 17 -111 25 -94
rect -25 -119 25 -111
<< polycont >>
rect -17 94 17 111
rect -17 -111 17 -94
<< locali >>
rect -105 145 -57 162
rect 57 145 105 162
rect -105 114 -88 145
rect 88 114 105 145
rect -25 94 -17 111
rect 17 94 25 111
rect -48 69 -31 77
rect -48 -77 -31 -69
rect 31 69 48 77
rect 31 -77 48 -69
rect -25 -111 -17 -94
rect 17 -111 25 -94
rect -105 -145 -88 -114
rect 88 -145 105 -114
rect -105 -162 -57 -145
rect 57 -162 105 -145
<< viali >>
rect -17 94 17 111
rect -48 -69 -31 69
rect 31 -69 48 69
rect -17 -111 17 -94
<< metal1 >>
rect -23 111 23 114
rect -23 94 -17 111
rect 17 94 23 111
rect -23 91 23 94
rect -51 69 -28 75
rect -51 -69 -48 69
rect -31 -69 -28 69
rect -51 -75 -28 -69
rect 28 69 51 75
rect 28 -69 31 69
rect 48 -69 51 69
rect 28 -75 51 -69
rect -23 -94 23 -91
rect -23 -111 -17 -94
rect 17 -111 23 -94
rect -23 -114 23 -111
<< properties >>
string FIXED_BBOX -96 -153 96 153
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.50 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
